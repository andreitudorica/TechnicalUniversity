---------------------------------------------------------------------------------------------------
--
-- Title       : \bcd-exces\
-- Design      : subiecte_2010
-- Author      : Andreea
-- Company     : a
--
---------------------------------------------------------------------------------------------------
--
-- File        : bcd-exces.vhd
-- Generated   : Sat May  7 18:41:14 2011
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {\bcd-exces\} architecture {\bcd-exces\}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity bcd-exces is
end bcd-exces;

--}} End of automatically maintained section

architecture bcd-exces3 of bcd-exces is
component bcd
	port 

	 -- enter your statements here --

end bcd-exces;
