-------------------------------------------------------------------------------
--
-- Title       : khkjhj
-- Design      : kjh
-- Author      : Ioana
-- Company     : UTCN
--
-------------------------------------------------------------------------------
--
-- File        : khkjhj.vhd
-- Generated   : Mon May 16 20:06:04 2011
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {khkjhj} architecture {khkjhj}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity khkjhj is
end khkjhj;

--}} End of automatically maintained section

architecture khkjhj of khkjhj is
begin

	 -- enter your statements here --

end khkjhj;
