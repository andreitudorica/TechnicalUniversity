--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:             12:22 PM, 4/15/99 *
--* Tested entity name:                        pr_sr_register *
--* File name contains tested entity: $DSN\src\serial_register.vhd *
--*************************************************************

library ieee;
use ieee.NUMERIC_STD.all;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity pr_sr_register_tb is
end pr_sr_register_tb;

architecture TB_ARCHITECTURE of pr_sr_register_tb is
	-- Component declaration of the tested unit
	component pr_sr_register
	port(
		nWRS : in std_logic;
		TXC : in std_logic;
		RESET : in std_logic;
		DATAS : in std_logic_vector(7 downto 0);
		INT : out std_logic;
		BUSY : out std_logic;
		TXD : out std_logic );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal nWRS : std_logic;
	signal TXC : std_logic;
	signal RESET : std_logic;
	signal DATAS : std_logic_vector(7 downto 0);
	-- Observed signals - signals mapped to the output ports of tested entity
	signal INT : std_logic;
	signal BUSY : std_logic;
	signal TXD : std_logic;

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : pr_sr_register
		port map
			(nWRS => nWRS,
			TXC => TXC,
			RESET => RESET,
			DATAS => DATAS,
			INT => INT,
			BUSY => BUSY,
			TXD => TXD );

	--Below VHDL code is an inserted .\compile\pr_sr.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	nWRS <= '1';
	TXC <= '1';
	DATAS <= "01010101";
	RESET <= '1';
    wait for 100 ns; --0 ps
	RESET <= '0';
    wait for 100 ns; --100 ns
	nWRS <= '0';
    wait for 100 ns; --200 ns
	nWRS <= '1';
    wait for 100 ns; --300 ns
	TXC <= '0';
    wait for 50 ns; --400 ns
	TXC <= '1';
    wait for 50 ns; --450 ns
	TXC <= '0';
    wait for 50 ns; --500 ns
	TXC <= '1';
    wait for 50 ns; --550 ns
	TXC <= '0';
    wait for 50 ns; --600 ns
	TXC <= '1';
    wait for 50 ns; --650 ns
	TXC <= '0';
    wait for 50 ns; --700 ns
	TXC <= '1';
    wait for 50 ns; --750 ns
	TXC <= '0';
    wait for 50 ns; --800 ns
	TXC <= '1';
    wait for 50 ns; --850 ns
	TXC <= '0';
    wait for 50 ns; --900 ns
	TXC <= '1';
    wait for 50 ns; --950 ns
	TXC <= '0';
    wait for 50 ns; --1 us
	TXC <= '1';
    wait for 50 ns; --1050 ns
	TXC <= '0';
    wait for 50 ns; --1100 ns
	TXC <= '1';
    wait for 150 ns; --1150 ns
	DATAS <= "10101010";
    wait for 100 ns; --1300 ns
	nWRS <= '0';
    wait for 100 ns; --1400 ns
	nWRS <= '1';
    wait for 100 ns; --1500 ns
	TXC <= '0';
    wait for 50 ns; --1600 ns
	TXC <= '1';
    wait for 50 ns; --1650 ns
	TXC <= '0';
    wait for 50 ns; --1700 ns
	TXC <= '1';
    wait for 50 ns; --1750 ns
	TXC <= '0';
    wait for 50 ns; --1800 ns
	TXC <= '1';
    wait for 50 ns; --1850 ns
	TXC <= '0';
    wait for 50 ns; --1900 ns
	TXC <= '1';
    wait for 50 ns; --1950 ns
	TXC <= '0';
    wait for 50 ns; --2 us
	TXC <= '1';
    wait for 50 ns; --2050 ns
	TXC <= '0';
    wait for 50 ns; --2100 ns
	TXC <= '1';
    wait for 50 ns; --2150 ns
	TXC <= '0';
    wait for 50 ns; --2200 ns
	TXC <= '1';
    wait for 50 ns; --2250 ns
	TXC <= '0';
    wait for 50 ns; --2300 ns
	TXC <= '1';
    wait for 150 ns; --2350 ns
	RESET <= '1';
    wait for 100 ns; --2500 ns
	RESET <= '0';
    wait for 100 ns; --2600 ns
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_pr_sr_register of pr_sr_register_tb is
	for TB_ARCHITECTURE
		for UUT : pr_sr_register
			use entity work.pr_sr_register(pr_sr_register);
		end for;
	end for;
end TESTBENCH_FOR_pr_sr_register;

