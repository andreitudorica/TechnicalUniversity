--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-HDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:               14:00, 99-05-20 *
--* Tested entity name:                              top_frqm *
--* File name contains tested entity: $DSN\compile\top_frqm.vhd *
--*************************************************************

library ieee;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity top_frqm_tb is
end top_frqm_tb;

architecture TB_ARCHITECTURE of top_frqm_tb is
	-- Component declaration of the tested unit
	component top_frqm
	port(
		F_INPUT : in std_logic;
		F_PATTERN : in std_logic;
		RESET : in std_logic;
		START : in std_logic;
		LED_A : out std_logic_vector(6 downto 0);
		LED_B : out std_logic_vector(6 downto 0);
		LED_C : out std_logic_vector(6 downto 0);
		LED_D : out std_logic_vector(6 downto 0) );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal F_INPUT : std_logic;
	signal F_PATTERN : std_logic;
	signal RESET : std_logic;
	signal START : std_logic;
	-- Observed signals - signals mapped to the output ports of tested entity
	signal LED_A : std_logic_vector(6 downto 0);
	signal LED_B : std_logic_vector(6 downto 0);
	signal LED_C : std_logic_vector(6 downto 0);
	signal LED_D : std_logic_vector(6 downto 0);

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : top_frqm
		port map
			(F_INPUT => F_INPUT,
			F_PATTERN => F_PATTERN,
			RESET => RESET,
			START => START,
			LED_A => LED_A,
			LED_B => LED_B,
			LED_C => LED_C,
			LED_D => LED_D );

	--Below VHDL code is an inserted .\compile\top_frqm.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	F_INPUT <= '0';
	F_PATTERN <= '0';
	RESET <= '1';
	START <= '0';
    wait for 50 ns; --0 ps
	F_INPUT <= '1';
    wait for 50 ns; --50 ns
	F_INPUT <= '0';
    wait for 50 ns; --100 ns
	F_INPUT <= '1';
    wait for 50 ns; --150 ns
	F_INPUT <= '0';
    wait for 50 ns; --200 ns
	F_INPUT <= '1';
    wait for 50 ns; --250 ns
	F_INPUT <= '0';
    wait for 50 ns; --300 ns
	F_INPUT <= '1';
    wait for 50 ns; --350 ns
	F_INPUT <= '0';
    wait for 50 ns; --400 ns
	F_INPUT <= '1';
    wait for 50 ns; --450 ns
	F_INPUT <= '0';
    wait for 50 ns; --500 ns
	F_INPUT <= '1';
    wait for 50 ns; --550 ns
	F_INPUT <= '0';
    wait for 50 ns; --600 ns
	F_INPUT <= '1';
    wait for 50 ns; --650 ns
	F_INPUT <= '0';
    wait for 50 ns; --700 ns
	F_INPUT <= '1';
    wait for 50 ns; --750 ns
	F_INPUT <= '0';
    wait for 50 ns; --800 ns
	F_INPUT <= '1';
    wait for 50 ns; --850 ns
	F_INPUT <= '0';
    wait for 50 ns; --900 ns
	F_INPUT <= '1';
    wait for 50 ns; --950 ns
	F_INPUT <= '0';
	F_PATTERN <= '1';
	RESET <= '0';
    wait for 50 ns; --1 us
	F_INPUT <= '1';
    wait for 50 ns; --1050 ns
	F_INPUT <= '0';
    wait for 50 ns; --1100 ns
	F_INPUT <= '1';
    wait for 50 ns; --1150 ns
	F_INPUT <= '0';
    wait for 50 ns; --1200 ns
	F_INPUT <= '1';
    wait for 50 ns; --1250 ns
	F_INPUT <= '0';
    wait for 50 ns; --1300 ns
	F_INPUT <= '1';
    wait for 50 ns; --1350 ns
	F_INPUT <= '0';
    wait for 50 ns; --1400 ns
	F_INPUT <= '1';
    wait for 50 ns; --1450 ns
	F_INPUT <= '0';
    wait for 50 ns; --1500 ns
	F_INPUT <= '1';
    wait for 50 ns; --1550 ns
	F_INPUT <= '0';
    wait for 50 ns; --1600 ns
	F_INPUT <= '1';
    wait for 50 ns; --1650 ns
	F_INPUT <= '0';
    wait for 50 ns; --1700 ns
	F_INPUT <= '1';
    wait for 50 ns; --1750 ns
	F_INPUT <= '0';
    wait for 50 ns; --1800 ns
	F_INPUT <= '1';
    wait for 50 ns; --1850 ns
	F_INPUT <= '0';
    wait for 50 ns; --1900 ns
	F_INPUT <= '1';
    wait for 50 ns; --1950 ns
	F_INPUT <= '0';
	F_PATTERN <= '0';
	START <= '1';
    wait for 50 ns; --2 us
	F_INPUT <= '1';
    wait for 50 ns; --2050 ns
	F_INPUT <= '0';
    wait for 50 ns; --2100 ns
	F_INPUT <= '1';
    wait for 50 ns; --2150 ns
	F_INPUT <= '0';
    wait for 50 ns; --2200 ns
	F_INPUT <= '1';
    wait for 50 ns; --2250 ns
	F_INPUT <= '0';
    wait for 50 ns; --2300 ns
	F_INPUT <= '1';
    wait for 50 ns; --2350 ns
	F_INPUT <= '0';
    wait for 50 ns; --2400 ns
	F_INPUT <= '1';
    wait for 50 ns; --2450 ns
	F_INPUT <= '0';
    wait for 50 ns; --2500 ns
	F_INPUT <= '1';
    wait for 50 ns; --2550 ns
	F_INPUT <= '0';
    wait for 50 ns; --2600 ns
	F_INPUT <= '1';
    wait for 50 ns; --2650 ns
	F_INPUT <= '0';
    wait for 50 ns; --2700 ns
	F_INPUT <= '1';
    wait for 50 ns; --2750 ns
	F_INPUT <= '0';
    wait for 50 ns; --2800 ns
	F_INPUT <= '1';
    wait for 50 ns; --2850 ns
	F_INPUT <= '0';
    wait for 50 ns; --2900 ns
	F_INPUT <= '1';
    wait for 50 ns; --2950 ns
	F_INPUT <= '0';
	F_PATTERN <= '1';
    wait for 50 ns; --3 us
	F_INPUT <= '1';
    wait for 50 ns; --3050 ns
	F_INPUT <= '0';
    wait for 50 ns; --3100 ns
	F_INPUT <= '1';
    wait for 50 ns; --3150 ns
	F_INPUT <= '0';
    wait for 50 ns; --3200 ns
	F_INPUT <= '1';
    wait for 50 ns; --3250 ns
	F_INPUT <= '0';
    wait for 50 ns; --3300 ns
	F_INPUT <= '1';
    wait for 50 ns; --3350 ns
	F_INPUT <= '0';
    wait for 50 ns; --3400 ns
	F_INPUT <= '1';
    wait for 50 ns; --3450 ns
	F_INPUT <= '0';
    wait for 50 ns; --3500 ns
	F_INPUT <= '1';
    wait for 50 ns; --3550 ns
	F_INPUT <= '0';
    wait for 50 ns; --3600 ns
	F_INPUT <= '1';
    wait for 50 ns; --3650 ns
	F_INPUT <= '0';
    wait for 50 ns; --3700 ns
	F_INPUT <= '1';
    wait for 50 ns; --3750 ns
	F_INPUT <= '0';
    wait for 50 ns; --3800 ns
	F_INPUT <= '1';
    wait for 50 ns; --3850 ns
	F_INPUT <= '0';
    wait for 50 ns; --3900 ns
	F_INPUT <= '1';
    wait for 50 ns; --3950 ns
	F_INPUT <= '0';
	F_PATTERN <= '0';
    wait for 50 ns; --4 us
	F_INPUT <= '1';
    wait for 50 ns; --4050 ns
	F_INPUT <= '0';
    wait for 50 ns; --4100 ns
	F_INPUT <= '1';
    wait for 50 ns; --4150 ns
	F_INPUT <= '0';
    wait for 50 ns; --4200 ns
	F_INPUT <= '1';
    wait for 50 ns; --4250 ns
	F_INPUT <= '0';
    wait for 50 ns; --4300 ns
	F_INPUT <= '1';
    wait for 50 ns; --4350 ns
	F_INPUT <= '0';
    wait for 50 ns; --4400 ns
	F_INPUT <= '1';
    wait for 50 ns; --4450 ns
	F_INPUT <= '0';
    wait for 50 ns; --4500 ns
	F_INPUT <= '1';
    wait for 50 ns; --4550 ns
	F_INPUT <= '0';
    wait for 50 ns; --4600 ns
	F_INPUT <= '1';
    wait for 50 ns; --4650 ns
	F_INPUT <= '0';
    wait for 50 ns; --4700 ns
	F_INPUT <= '1';
    wait for 50 ns; --4750 ns
	F_INPUT <= '0';
    wait for 50 ns; --4800 ns
	F_INPUT <= '1';
    wait for 50 ns; --4850 ns
	F_INPUT <= '0';
    wait for 50 ns; --4900 ns
	F_INPUT <= '1';
    wait for 50 ns; --4950 ns
	F_INPUT <= '0';
	F_PATTERN <= '1';
    wait for 50 ns; --5 us
	F_INPUT <= '1';
    wait for 50 ns; --5050 ns
	F_INPUT <= '0';
    wait for 50 ns; --5100 ns
	F_INPUT <= '1';
    wait for 50 ns; --5150 ns
	F_INPUT <= '0';
    wait for 50 ns; --5200 ns
	F_INPUT <= '1';
    wait for 50 ns; --5250 ns
	F_INPUT <= '0';
    wait for 50 ns; --5300 ns
	F_INPUT <= '1';
    wait for 50 ns; --5350 ns
	F_INPUT <= '0';
    wait for 50 ns; --5400 ns
	F_INPUT <= '1';
    wait for 50 ns; --5450 ns
	F_INPUT <= '0';
    wait for 50 ns; --5500 ns
	F_INPUT <= '1';
    wait for 50 ns; --5550 ns
	F_INPUT <= '0';
    wait for 50 ns; --5600 ns
	F_INPUT <= '1';
    wait for 50 ns; --5650 ns
	F_INPUT <= '0';
    wait for 50 ns; --5700 ns
	F_INPUT <= '1';
    wait for 50 ns; --5750 ns
	F_INPUT <= '0';
    wait for 50 ns; --5800 ns
	F_INPUT <= '1';
    wait for 50 ns; --5850 ns
	F_INPUT <= '0';
    wait for 50 ns; --5900 ns
	F_INPUT <= '1';
    wait for 50 ns; --5950 ns
	F_INPUT <= '0';
	F_PATTERN <= '0';
    wait for 50 ns; --6 us
	F_INPUT <= '1';
    wait for 50 ns; --6050 ns
	F_INPUT <= '0';
    wait for 50 ns; --6100 ns
	F_INPUT <= '1';
    wait for 50 ns; --6150 ns
	F_INPUT <= '0';
    wait for 50 ns; --6200 ns
	F_INPUT <= '1';
    wait for 50 ns; --6250 ns
	F_INPUT <= '0';
    wait for 50 ns; --6300 ns
	F_INPUT <= '1';
    wait for 50 ns; --6350 ns
	F_INPUT <= '0';
    wait for 50 ns; --6400 ns
	F_INPUT <= '1';
	START <= '0';
    wait for 50 ns; --6450 ns
	F_INPUT <= '0';
    wait for 50 ns; --6500 ns
	F_INPUT <= '1';
    wait for 50 ns; --6550 ns
	F_INPUT <= '0';
    wait for 50 ns; --6600 ns
	F_INPUT <= '1';
    wait for 50 ns; --6650 ns
	F_INPUT <= '0';
    wait for 50 ns; --6700 ns
	F_INPUT <= '1';
    wait for 50 ns; --6750 ns
	F_INPUT <= '0';
    wait for 50 ns; --6800 ns
	F_INPUT <= '1';
    wait for 50 ns; --6850 ns
	F_INPUT <= '0';
    wait for 50 ns; --6900 ns
	F_INPUT <= '1';
    wait for 50 ns; --6950 ns
	F_INPUT <= '0';
	F_PATTERN <= '1';
    wait for 50 ns; --7 us
	F_INPUT <= '1';
    wait for 50 ns; --7050 ns
	F_INPUT <= '0';
    wait for 50 ns; --7100 ns
	F_INPUT <= '1';
    wait for 50 ns; --7150 ns
	F_INPUT <= '0';
    wait for 50 ns; --7200 ns
	F_INPUT <= '1';
    wait for 50 ns; --7250 ns
	F_INPUT <= '0';
    wait for 50 ns; --7300 ns
	F_INPUT <= '1';
    wait for 50 ns; --7350 ns
	F_INPUT <= '0';
    wait for 50 ns; --7400 ns
	F_INPUT <= '1';
    wait for 50 ns; --7450 ns
	F_INPUT <= '0';
    wait for 50 ns; --7500 ns
	F_INPUT <= '1';
    wait for 50 ns; --7550 ns
	F_INPUT <= '0';
    wait for 50 ns; --7600 ns
	F_INPUT <= '1';
    wait for 50 ns; --7650 ns
	F_INPUT <= '0';
    wait for 50 ns; --7700 ns
	F_INPUT <= '1';
    wait for 50 ns; --7750 ns
	F_INPUT <= '0';
    wait for 50 ns; --7800 ns
	F_INPUT <= '1';
    wait for 50 ns; --7850 ns
	F_INPUT <= '0';
    wait for 50 ns; --7900 ns
	F_INPUT <= '1';
    wait for 50 ns; --7950 ns
	F_INPUT <= '0';
    wait for 1 ps; --8 us
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_top_frqm of top_frqm_tb is
	for TB_ARCHITECTURE
		for UUT : top_frqm
			use entity work.top_frqm(top_frqm);
		end for;
	end for;
end TESTBENCH_FOR_top_frqm;

