--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:               4:12 PM, 4/7/99 *
--* Tested entity name:                                   ram *
--* File name contains tested entity:        $DSN\src\ram.vhd *
--*************************************************************

library ieee;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity ram_tb is
	-- Generic declarations of the tested unit
	generic(
		AddSize : INTEGER := 4 );
end ram_tb;

architecture TB_ARCHITECTURE of ram_tb is
	-- Component declaration of the tested unit
	component ram
	generic(
		AddSize : INTEGER := 4 );
	port(
		nRD : in std_logic;
		nWR : in std_logic;
		nCS : in std_logic;
		DATA : inout std_logic_vector(7 downto 0);
		ADDRESS : in std_logic_vector((AddSize-1) downto 0) );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal nRD : std_logic;
	signal nWR : std_logic;
	signal nCS : std_logic;
	signal DATA : std_logic_vector(7 downto 0);
	signal ADDRESS : std_logic_vector((AddSize-1) downto 0);
	-- Observed signals - signals mapped to the output ports of tested entity

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : ram
		port map
			(nRD => nRD,
			nWR => nWR,
			nCS => nCS,
			DATA => DATA,
			ADDRESS => ADDRESS );

	--Below VHDL code is an inserted .\compile\ram.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	nWR <= '1';
	ADDRESS <= "0000";
	nRD <= '1';
	nCS <= '0';
	DATA <= "00000000";
    wait for 100 ns; --0 ps
	nWR <= '0';
    wait for 100 ns; --100 ns
	nWR <= '1';
    wait for 100 ns; --200 ns
	ADDRESS <= "0001";
	DATA <= "00000001";
    wait for 100 ns; --300 ns
	nWR <= '0';
    wait for 100 ns; --400 ns
	nWR <= '1';
    wait for 100 ns; --500 ns
	ADDRESS <= "0010";
	DATA <= "00000010";
    wait for 100 ns; --600 ns
	nWR <= '0';
    wait for 100 ns; --700 ns
	nWR <= '1';
    wait for 100 ns; --800 ns
	ADDRESS <= "0011";
	DATA <= "00000011";
    wait for 100 ns; --900 ns
	nWR <= '0';
    wait for 100 ns; --1 us
	nWR <= '1';
    wait for 100 ns; --1100 ns
	ADDRESS <= "0100";
	DATA <= "00000100";
    wait for 100 ns; --1200 ns
	nWR <= '0';
    wait for 100 ns; --1300 ns
	nWR <= '1';
    wait for 100 ns; --1400 ns
	ADDRESS <= "0101";
	DATA <= "00000101";
    wait for 100 ns; --1500 ns
	nWR <= '0';
    wait for 100 ns; --1600 ns
	nWR <= '1';
    wait for 100 ns; --1700 ns
	ADDRESS <= "0110";
	DATA <= "00000110";
    wait for 100 ns; --1800 ns
	nWR <= '0';
    wait for 100 ns; --1900 ns
	nWR <= '1';
    wait for 100 ns; --2 us
	ADDRESS <= "0111";
	DATA <= "00000111";
    wait for 100 ns; --2100 ns
	nWR <= '0';
    wait for 100 ns; --2200 ns
	nWR <= '1';
    wait for 100 ns; --2300 ns
	ADDRESS <= "0000";
	DATA <= "ZZZZZZZZ";
    wait for 100 ns; --2400 ns
	nRD <= '0';
    wait for 100 ns; --2500 ns
	nRD <= '1';
    wait for 100 ns; --2600 ns
	ADDRESS <= "0001";
    wait for 100 ns; --2700 ns
	nRD <= '0';
    wait for 100 ns; --2800 ns
	nRD <= '1';
    wait for 100 ns; --2900 ns
	ADDRESS <= "0010";
    wait for 100 ns; --3 us
	nRD <= '0';
    wait for 100 ns; --3100 ns
	nRD <= '1';
    wait for 100 ns; --3200 ns
	ADDRESS <= "0011";
    wait for 100 ns; --3300 ns
	nRD <= '0';
    wait for 100 ns; --3400 ns
	nRD <= '1';
	DATA <= "ZZZZZZZZ";
    wait for 100 ns; --3500 ns
	ADDRESS <= "0100";
    wait for 100 ns; --3600 ns
	nRD <= '0';
    wait for 100 ns; --3700 ns
	nRD <= '1';
    wait for 100 ns; --3800 ns
	ADDRESS <= "0101";
    wait for 100 ns; --3900 ns
	nRD <= '0';
    wait for 100 ns; --4 us
	nRD <= '1';
    wait for 100 ns; --4100 ns
	ADDRESS <= "0110";
    wait for 100 ns; --4200 ns
	nRD <= '0';
    wait for 100 ns; --4300 ns
	nRD <= '1';
    wait for 100 ns; --4400 ns
	ADDRESS <= "0111";
    wait for 100 ns; --4500 ns
	nRD <= '0';
    wait for 100 ns; --4600 ns
	nRD <= '1';
    wait for 100 ns; --4700 ns
	ADDRESS <= "1000";
    wait for 100 ns; --4800 ns
	nRD <= '0';
	wait for 100 ns; --4900 ns
	nRD <= '1';
	wait for 100 ns; --5 us
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_ram of ram_tb is
	for TB_ARCHITECTURE
		for UUT : ram
			use entity work.ram(ram);
		end for;
	end for;
end TESTBENCH_FOR_ram;

