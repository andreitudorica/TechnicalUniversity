entity ROM is
	port(I: in natural;
	     Y: out bit_vector(0 to 15));
end ROM;

architecture arh_ROM of ROM is
begin
	process(I)
	type ROM is array(0 to 15) of bit_vector(0 to 15); --????
	variable X:ROM;
	begin		   
		X(0) :="1000000000000000";
		X(1) :="0100000000000000";
		X(2) :="0010000000000000";
		X(3) :="0001000000000000";
		X(4) :="0000100000000000";
		X(5) :="0000010000000000";
		X(6) :="0000001000000000";
		X(7) :="0000000100000000";
		X(8) :="0000000010000000";
		X(9) :="0000000001000000";
		X(10):="0000000000100000";
		X(11):="0000000000010000";
		X(12):="0000000000001000";
		X(13):="0000000000000100";
		X(14):="0000000000000010";
		X(15):="0000000000000001";
		
		Y<=X(I);
	end process;
end arh_ROM;